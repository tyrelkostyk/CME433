module parity_conventional( D, F );

input [6:0] D;
output F;

assign F = (~D[0] & D[1] & ~D[2] & D[3] & D[5]) ^
        (D[2] & ~D[3] & D[5]) ^
        (D[0] & ~D[1] & ~D[2] & ~D[3] & ~D[4] & ~D[6]) ^
        (D[0] & D[1] & D[2] & ~D[3] & D[5]) ^
        (D[0] & ~D[1] & ~D[3]) ^ 
        (~D[0] & D[1] & D[3] & D[5] & ~D[6]) ^ 
        (~D[0] & D[2] & D[3] & D[5] & ~D[6]) ^ 
        (~D[0] & D[1] & D[2] & ~D[3] & ~D[4] & ~D[5] & D[6]) ^ 
        (~D[0] & D[2]) ^ 
        (~D[0] & D[1] & ~D[2] & ~D[6]) ^ 
        (~D[1] & ~D[2] & ~D[3] & ~D[4]);

endmodule
